ADDED NEW CONTENT